module screenbuffer(
	input wire wren;
	input wire [7:0] address_a;
	wire [7:0]
);